module top_module( output one );

// Insert your code here
    assign one = 2'b01;
endmodule